module top_module # (
    parameter N = 16,      // Number of bits input
    parameter NUM_FIRS = 8, // Number of FIR filters

    parameter DELAYS = 62, 

    parameter GAIN_1 = 2, 
    parameter GAIN_2 = 4,
    parameter GAIN_3 = 6,
    parameter GAIN_4 = 8,
    parameter GAIN_5 = 10,
    parameter GAIN_6 = 12,
    parameter GAIN_7 = 14,
    parameter GAIN_8 = 16       


) (
    input  clk,
    input  rst,
    input  ena,
    input  signed [N-1:0] x_in,
    
    output reg signed [N*2-1:0] y_out_1,
    output reg signed [N*2-1:0] y_out_2,
    output reg signed [N*2-1:0] y_out_3,
    output reg signed [N*2-1:0] y_out_4,
    output reg signed [N*2-1:0] y_out_5,
    output reg signed [N*2-1:0] y_out_6,
    output reg signed [N*2-1:0] y_out_7,
    output reg signed [N*2-1:0] y_out_8,
    output reg signed [N*2-1:0] y_out
);

    wire [N*2-1:0] y_out_1_to_gain;
    wire [N*2-1:0] y_out_2_to_gain;
    wire [N*2-1:0] y_out_3_to_gain;
    wire [N*2-1:0] y_out_4_to_gain;
    wire [N*2-1:0] y_out_5_to_gain;
    wire [N*2-1:0] y_out_6_to_gain;
    wire [N*2-1:0] y_out_7_to_gain;
    wire [N*2-1:0] y_out_8_to_gain;
   
	//parameter INTEGER_COEFF_WIDTH = 6; // Width of each coefficient in bits
    // parameter logic [5:0] DELAYS [1:8] = { // Use array have 8 elements , each element have 6bits
    //     6'd62, 
    //     6'd42,
    //     6'd48,
    //     6'd48,
    //     6'd48,
    //     6'd50,
    //     6'd52,
    //     6'd52      
    // };

   // parameter [(52+1)*N-1:0] COEFFICIENTS [1:8]

    // parameter [NUM_FIRS*64-1:0] DELAYS = '{3, 4, 5, 6, 7, 8, 9, 10}; // Array of DELAYS for each FIR filter
    // parameter [NUM_FIRS-1:0] COEFFICIENTS = '{32'h12345678, 32'h23456789, 32'h3456789A, 32'h456789AB, 32'h56789ABC, 32'h6789ABCD, 32'h789ABCDE, 32'h89ABCDEF}; // Array of coefficients for each FIR filter
    parameter [(DELAYS+1)*8-1:0] b_1 = {
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111110,
        8'b11111110,
        8'b11111110,
        8'b11111111,
        8'b0,
        8'b1,
        8'b10,
        8'b100,
        8'b101,
        8'b101,
        8'b101,
        8'b11,
        8'b11111111,
        8'b11111011,
        8'b11110110,
        8'b11110001,
        8'b11101101,
        8'b11101100,
        8'b11101110,
        8'b11110100,
        8'b0,
        8'b1111,
        8'b100010,
        8'b110111,
        8'b1001100,
        8'b1100000,
        8'b1101111,
        8'b1111001,
        8'b1111101,
        8'b1111001,
        8'b1101111,
        8'b1100000,
        8'b1001100,
        8'b110111,
        8'b100010,
        8'b1111,
        8'b0,
        8'b11110100,
        8'b11101110,
        8'b11101100,
        8'b11101101,
        8'b11110001,
        8'b11110110,
        8'b11111011,
        8'b11111111,
        8'b11,
        8'b101,
        8'b101,
        8'b101,
        8'b100,
        8'b10,
        8'b1,
        8'b0,
        8'b11111111,
        8'b11111110,
        8'b11111110,
        8'b11111110,
        8'b11111111,
        8'b11111111,
        8'b11111111
    };

    parameter [(DELAYS+1)*N-1:0] b_2 = {
        8'b11111111,
        8'b11111111,
        8'b0,
        8'b1,
        8'b10,
        8'b10,
        8'b10,
        8'b11111111,
        8'b11111100,
        8'b11111001,
        8'b11111000,
        8'b11111010,
        8'b11111110,
        8'b10,
        8'b10,
        8'b11111111,
        8'b11111100,
        8'b11111011,
        8'b11,
        8'b10010,
        8'b100010,
        8'b101010,
        8'b11111,
        8'b11111111,
        8'b11010100,
        8'b10101101,
        8'b10011110,
        8'b10110011,
        8'b11101001,
        8'b101101,
        8'b1100110,
        8'b1111100,
        8'b1100110,
        8'b101101,
        8'b11101001,
        8'b10110011,
        8'b10011110,
        8'b10101101,
        8'b11010100,
        8'b11111111,
        8'b11111,
        8'b101010,
        8'b100010,
        8'b10010,
        8'b11,
        8'b11111011,
        8'b11111100,
        8'b11111111,
        8'b10,
        8'b10,
        8'b11111110,
        8'b11111010,
        8'b11111000,
        8'b11111001,
        8'b11111100,
        8'b11111111,
        8'b10,
        8'b10,
        8'b10,
        8'b1,
        8'b0,
        8'b11111111,
        8'b11111111
    };

    parameter [(DELAYS+1)*N-1:0] b_3 = {
        8'b11111111,
        8'b00000000,
        8'b00000001,
        8'b00000001,
        8'b11111111,
        8'b11111101,
        8'b11111100,
        8'b00000000,
        8'b00000101,
        8'b00000110,
        8'b00000001,
        8'b11111010,
        8'b11111001,
        8'b11111101,
        8'b00000001,
        8'b11111111,
        8'b11111101,
        8'b00000100,
        8'b00010001,
        8'b00010010,
        8'b11111001,
        8'b11010101,
        8'b11010000,
        8'b00000000,
        8'b01000001,
        8'b01010010,
        8'b00010011,
        8'b10110011,
        8'b10001111,
        8'b11010001,
        8'b01000100,
        8'b01111100,
        8'b01000100,
        8'b11010001,
        8'b10001111,
        8'b10110011,
        8'b00010011,
        8'b01010010,
        8'b01000001,
        8'b00000000,
        8'b11010000,
        8'b11010101,
        8'b11111001,
        8'b00010010,
        8'b00010001,
        8'b00000100,
        8'b11111101,
        8'b11111111,
        8'b00000001,
        8'b11111101,
        8'b11111001,
        8'b11111010,
        8'b00000001,
        8'b00000110,
        8'b00000101,
        8'b00000000,
        8'b11111100,
        8'b11111101,
        8'b11111111,
        8'b00000001,
        8'b00000001,
        8'b00000000,
        8'b11111111
    };

    parameter [(DELAYS+1)*N-1:0] b_4 = {
        8'b11111111,
        8'b00000000,
        8'b00000000,
        8'b11111110,
        8'b11111110,
        8'b00000001,
        8'b00000011,
        8'b11111111,
        8'b11111010,
        8'b11111101,
        8'b00000110,
        8'b00000101,
        8'b11111100,
        8'b11111010,
        8'b00000000,
        8'b11111111,
        8'b11111111,
        8'b00001001,
        8'b00001001,
        8'b11101101,
        8'b11100010,
        8'b00010001,
        8'b00110111,
        8'b11111111,
        8'b10110010,
        8'b11011101,
        8'b01010010,
        8'b01001100,
        8'b11000000,
        8'b10010000,
        8'b00011000,
        8'b01111100,
        8'b00011000,
        8'b10010000,
        8'b11000000,
        8'b01001100,
        8'b01010010,
        8'b11011101,
        8'b10110010,
        8'b11111111,
        8'b00110111,
        8'b00010001,
        8'b11100010,
        8'b11101101,
        8'b00001001,
        8'b00001001,
        8'b11111111,
        8'b11111111,
        8'b00000000,
        8'b11111010,
        8'b11111100,
        8'b00000101,
        8'b00000110,
        8'b11111101,
        8'b11111010,
        8'b11111111,
        8'b00000011,
        8'b00000001,
        8'b11111110,
        8'b11111110,
        8'b00000000,
        8'b00000000,
        8'b11111111
    };

    parameter [(DELAYS+1)*N-1:0] b_5 = {
        8'b00000000,
        8'b00000000,
        8'b11111111,
        8'b11111110,
        8'b00000001,
        8'b00000001,
        8'b11111100,
        8'b00000000,
        8'b00000101,
        8'b11111101,
        8'b11111001,
        8'b00000101,
        8'b00000011,
        8'b11111010,
        8'b11111111,
        8'b11111111,
        8'b00000000,
        8'b00001001,
        8'b11110110,
        8'b11101101,
        8'b00011101,
        8'b00010001,
        8'b11001000,
        8'b00000000,
        8'b01001101,
        8'b11011101,
        8'b10101101,
        8'b01001100,
        8'b00111111,
        8'b10010000,
        8'b11100111,
        8'b01111100,
        8'b11100111,
        8'b10010000,
        8'b00111111,
        8'b01001100,
        8'b10101101,
        8'b11011101,
        8'b01001101,
        8'b00000000,
        8'b11001000,
        8'b00010001,
        8'b00011101,
        8'b11101101,
        8'b11110110,
        8'b00001001,
        8'b00000000,
        8'b11111111,
        8'b11111111,
        8'b11111010,
        8'b00000011,
        8'b00000101,
        8'b11111001,
        8'b11111101,
        8'b00000101,
        8'b00000000,
        8'b11111100,
        8'b00000001,
        8'b00000001,
        8'b11111110,
        8'b11111111,
        8'b00000000,
        8'b00000000
    };

    parameter [(DELAYS+1)*N-1:0] b_6 = {
        8'b00000000,
        8'b00000000,
        8'b11111110,
        8'b00000001,
        8'b00000000,
        8'b11111101,
        8'b00000011,
        8'b11111111,
        8'b11111010,
        8'b00000110,
        8'b11111110,
        8'b11111010,
        8'b00000110,
        8'b11111101,
        8'b11111110,
        8'b11111111,
        8'b00000010,
        8'b00000100,
        8'b11101110,
        8'b00010010,
        8'b00000110,
        8'b11010101,
        8'b00101111,
        8'b11111111,
        8'b10111110,
        8'b01010010,
        8'b11101100,
        8'b10110011,
        8'b01110000,
        8'b11010001,
        8'b10111011,
        8'b01111100,
        8'b10111011,
        8'b11010001,
        8'b01110000,
        8'b10110011,
        8'b11101100,
        8'b01010010,
        8'b10111110,
        8'b11111111,
        8'b00101111,
        8'b11010101,
        8'b00000110,
        8'b00010010,
        8'b11101110,
        8'b00000100,
        8'b00000010,
        8'b11111111,
        8'b11111110,
        8'b11111101,
        8'b00000110,
        8'b11111010,
        8'b11111110,
        8'b00000110,
        8'b11111010,
        8'b11111111,
        8'b00000011,
        8'b11111101,
        8'b00000000,
        8'b00000001,
        8'b11111110,
        8'b00000000,
        8'b00000000
    };

    parameter [(DELAYS+1)*N-1:0] b_7 = {
        8'b00000000,
        8'b11111111,
        8'b11111111,
        8'b00000001,
        8'b11111101,
        8'b00000010,
        8'b11111101,
        8'b00000000,
        8'b00000011,
        8'b11111001,
        8'b00000111,
        8'b11111010,
        8'b00000001,
        8'b00000010,
        8'b11111101,
        8'b11111111,
        8'b00000011,
        8'b11111011,
        8'b11111100,
        8'b00010010,
        8'b11011101,
        8'b00101010,
        8'b11100000,
        8'b00000000,
        8'b00101011,
        8'b10101101,
        8'b01100001,
        8'b10110011,
        8'b00010110,
        8'b00101101,
        8'b10011001,
        8'b01111100,
        8'b10011001,
        8'b00101101,
        8'b00010110,
        8'b10110011,
        8'b01100001,
        8'b10101101,
        8'b00101011,
        8'b00000000,
        8'b11100000,
        8'b00101010,
        8'b11011101,
        8'b00010010,
        8'b11111100,
        8'b11111011,
        8'b00000011,
        8'b11111111,
        8'b11111101,
        8'b00000010,
        8'b00000001,
        8'b11111010,
        8'b00000111,
        8'b11111001,
        8'b00000011,
        8'b00000000,
        8'b11111101,
        8'b00000010,
        8'b11111101,
        8'b00000001,
        8'b11111111,
        8'b11111111,
        8'b00000000
    };

    parameter [(DELAYS+1)*N-1:0] b_8 = {
        8'b00000000,
        8'b11111111,
        8'b00000000,
        8'b11111110,
        8'b00000001,
        8'b11111110,
        8'b00000000,
        8'b11111111,
        8'b11111110,
        8'b00000010,
        8'b11111011,
        8'b00000101,
        8'b11111010,
        8'b00000101,
        8'b11111100,
        8'b11111111,
        8'b00000100,
        8'b11110110,
        8'b00001110,
        8'b11101101,
        8'b00010011,
        8'b11101110,
        8'b00001011,
        8'b11111111,
        8'b11110000,
        8'b00100010,
        8'b11001000,
        8'b01001100,
        8'b10011111,
        8'b01101111,
        8'b10000110,
        8'b01111101,
        8'b10000110,
        8'b01101111,
        8'b10011111,
        8'b01001100,
        8'b11001000,
        8'b00100010,
        8'b11110000,
        8'b11111111,
        8'b00001011,
        8'b11101110,
        8'b00010011,
        8'b11101101,
        8'b00001110,
        8'b11110110,
        8'b00000100,
        8'b11111111,
        8'b11111100,
        8'b00000101,
        8'b11111010,
        8'b00000101,
        8'b11111011,
        8'b00000010,
        8'b11111110,
        8'b11111111,
        8'b00000000,
        8'b11111110,
        8'b00000001,
        8'b11111110,
        8'b00000000,
        8'b11111111,
        8'b00000000
    };

    fir_n #(.DELAYS(DELAYS), 
            .N(N)) fir_1 (
        .clk(clk), 
        .rst(rst), 
        .ena(ena), 
        .b(b_1), 
        .x_in(x_in), 
        .y_out(y_out_1_to_gain)
    );

    fir_n #(.DELAYS(DELAYS), 
            .N(N)) fir_2 (
        .clk(clk), 
        .rst(rst), 
        .ena(ena), 
        .b(b_2), 
        .x_in(x_in), 
        .y_out(y_out_2_to_gain)
    );

    fir_n #(.DELAYS(DELAYS), 
            .N(N)) fir_3 (
        .clk(clk), 
        .rst(rst), 
        .ena(ena), 
        .b(b_3), 
        .x_in(x_in), 
        .y_out(y_out_3_to_gain)
    );

    fir_n #(.DELAYS(DELAYS), 
            .N(N)) fir_4 (
        .clk(clk), 
        .rst(rst), 
        .ena(ena), 
        .b(b_4), 
        .x_in(x_in), 
        .y_out(y_out_4_to_gain)
    );

    fir_n #(.DELAYS(DELAYS), 
            .N(N)) fir_5 (
        .clk(clk), 
        .rst(rst), 
        .ena(ena), 
        .b(b_5), 
        .x_in(x_in), 
        .y_out(y_out_5_to_gain)
    );

    fir_n #(.DELAYS(DELAYS), 
            .N(N)) fir_6 (
        .clk(clk), 
        .rst(rst), 
        .ena(ena), 
        .b(b_6), 
        .x_in(x_in), 
        .y_out(y_out_6_to_gain)
    );

    fir_n #(.DELAYS(DELAYS), 
            .N(N)) fir_7 (
        .clk(clk), 
        .rst(rst), 
        .ena(ena), 
        .b(b_7), 
        .x_in(x_in), 
        .y_out(y_out_7_to_gain)
    );

    fir_n #(.DELAYS(DELAYS),
            .N(N)) fir_8 (
        .clk(clk), 
        .rst(rst), 
        .ena(ena), 
        .b(b_8), 
        .x_in(x_in), 
        .y_out(y_out_8_to_gain)
    );

	always@(posedge clk or negedge rst) begin
		if(~rst) begin
             y_out_1 <= 0;
             y_out_2 <= 0;
             y_out_3 <= 0;
             y_out_4 <= 0;
             y_out_5 <= 0;
             y_out_6 <= 0;
             y_out_7 <= 0;
             y_out_8 <= 0;
             y_out <= 0;

		end else if(ena) begin
			 y_out_1 <=y_out_1_to_gain * GAIN_1;
             y_out_2 <=y_out_2_to_gain * GAIN_2;
             y_out_3 <=y_out_3_to_gain * GAIN_3;
             y_out_4 <=y_out_4_to_gain * GAIN_4;
             y_out_5 <=y_out_5_to_gain * GAIN_5;
             y_out_6 <=y_out_6_to_gain * GAIN_6;
             y_out_7 <=y_out_7_to_gain * GAIN_7;
             y_out_8 <=y_out_8_to_gain * GAIN_8;
             y_out <= y_out_1 + y_out_2 + y_out_3 + y_out_4 + y_out_5 + y_out_6 + y_out_7 + y_out_8;
		end
	end

endmodule