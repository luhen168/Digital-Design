module cnt_y_thousand_hundred (
    input clk,
    input rst,
    input pulse_increase, pulse_decrease, enable_cnt_y,
    output [6:0] cnt_y_thousand_hundred // var type net is wire 
);

    reg [6:0] cnt;
    reg pre_increase, pre_decrease; 

    always @(posedge clk or negedge rst) begin
        if (~rst) begin
            cnt <= 7'd0;
            pre_increase <= 1;
            pre_decrease <= 1; 
        end else begin
            if (enable_cnt_y) begin
                if(pulse_increase != pre_increase) begin
                    pre_increase <= pulse_increase;
                    if(pulse_increase == 0) begin 
                        if (cnt == 7'd99) cnt <= 7'd0;
                        else cnt <= cnt + 1;
                    end
                end else if (pulse_decrease != pre_decrease) begin
                    pre_decrease <= pulse_decrease;
                    if(pulse_decrease) begin
                        if (cnt == 7'd00) cnt <= 7'd99;
                        else cnt <= cnt - 1;
                    end
                end
            end 
        end
    end
    assign cnt_y_thousand_hundred = cnt;
endmodule