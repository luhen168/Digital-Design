module top_7_seg(
	input [13:0]  bin,
	output [13:0]  display
);

	assign display [6:0] =  bin[6:0];
	assign display [13:7] = bin[13:7];
endmodule 	